module phase1_tb ();

phase1 dut (.*);