module phase1 (
    ports
);

    
endmodule